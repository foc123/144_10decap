*-- interposer PDN spice model 'interposer1' for AC analysis
*-- Total unit cell #: 81 (9x9)

.param cellno=81
.param r_int_cell='1e-3'
.param l_int_cell='1e-10'
.param c_int_cell='1e-11'

xdint_0_0 ndint_x_0_0 ndint_x_1000_0 ndint_y_0_0 ndint_y_0_1000 ndint_xy_0_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_1 ndint_x_1000_0 ndint_x_2000_0 ndint_y_1000_0 ndint_y_1000_1000 ndint_xy_1000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_2 ndint_x_2000_0 ndint_x_3000_0 ndint_y_2000_0 ndint_y_2000_1000 ndint_xy_2000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_3 ndint_x_3000_0 ndint_x_4000_0 ndint_y_3000_0 ndint_y_3000_1000 ndint_xy_3000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_4 ndint_x_4000_0 ndint_x_5000_0 ndint_y_4000_0 ndint_y_4000_1000 ndint_xy_4000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_5 ndint_x_5000_0 ndint_x_6000_0 ndint_y_5000_0 ndint_y_5000_1000 ndint_xy_5000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_6 ndint_x_6000_0 ndint_x_7000_0 ndint_y_6000_0 ndint_y_6000_1000 ndint_xy_6000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_7 ndint_x_7000_0 ndint_x_8000_0 ndint_y_7000_0 ndint_y_7000_1000 ndint_xy_7000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_0_8 ndint_x_8000_0 ndint_x_9000_0 ndint_y_8000_0 ndint_y_8000_1000 ndint_xy_8000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_0 ndint_x_0_1000 ndint_x_1000_1000 ndint_y_0_1000 ndint_y_0_2000 ndint_xy_0_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_1 ndint_x_1000_1000 ndint_x_2000_1000 ndint_y_1000_1000 ndint_y_1000_2000 ndint_xy_1000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_2 ndint_x_2000_1000 ndint_x_3000_1000 ndint_y_2000_1000 ndint_y_2000_2000 ndint_xy_2000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_3 ndint_x_3000_1000 ndint_x_4000_1000 ndint_y_3000_1000 ndint_y_3000_2000 ndint_xy_3000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_4 ndint_x_4000_1000 ndint_x_5000_1000 ndint_y_4000_1000 ndint_y_4000_2000 ndint_xy_4000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_5 ndint_x_5000_1000 ndint_x_6000_1000 ndint_y_5000_1000 ndint_y_5000_2000 ndint_xy_5000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_6 ndint_x_6000_1000 ndint_x_7000_1000 ndint_y_6000_1000 ndint_y_6000_2000 ndint_xy_6000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_7 ndint_x_7000_1000 ndint_x_8000_1000 ndint_y_7000_1000 ndint_y_7000_2000 ndint_xy_7000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_1_8 ndint_x_8000_1000 ndint_x_9000_1000 ndint_y_8000_1000 ndint_y_8000_2000 ndint_xy_8000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_0 ndint_x_0_2000 ndint_x_1000_2000 ndint_y_0_2000 ndint_y_0_3000 ndint_xy_0_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_1 ndint_x_1000_2000 ndint_x_2000_2000 ndint_y_1000_2000 ndint_y_1000_3000 ndint_xy_1000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_2 ndint_x_2000_2000 ndint_x_3000_2000 ndint_y_2000_2000 ndint_y_2000_3000 ndint_xy_2000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_3 ndint_x_3000_2000 ndint_x_4000_2000 ndint_y_3000_2000 ndint_y_3000_3000 ndint_xy_3000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_4 ndint_x_4000_2000 ndint_x_5000_2000 ndint_y_4000_2000 ndint_y_4000_3000 ndint_xy_4000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_5 ndint_x_5000_2000 ndint_x_6000_2000 ndint_y_5000_2000 ndint_y_5000_3000 ndint_xy_5000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_6 ndint_x_6000_2000 ndint_x_7000_2000 ndint_y_6000_2000 ndint_y_6000_3000 ndint_xy_6000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_7 ndint_x_7000_2000 ndint_x_8000_2000 ndint_y_7000_2000 ndint_y_7000_3000 ndint_xy_7000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_2_8 ndint_x_8000_2000 ndint_x_9000_2000 ndint_y_8000_2000 ndint_y_8000_3000 ndint_xy_8000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_0 ndint_x_0_3000 ndint_x_1000_3000 ndint_y_0_3000 ndint_y_0_4000 ndint_xy_0_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_1 ndint_x_1000_3000 ndint_x_2000_3000 ndint_y_1000_3000 ndint_y_1000_4000 ndint_xy_1000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_2 ndint_x_2000_3000 ndint_x_3000_3000 ndint_y_2000_3000 ndint_y_2000_4000 ndint_xy_2000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_3 ndint_x_3000_3000 ndint_x_4000_3000 ndint_y_3000_3000 ndint_y_3000_4000 ndint_xy_3000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_4 ndint_x_4000_3000 ndint_x_5000_3000 ndint_y_4000_3000 ndint_y_4000_4000 ndint_xy_4000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_5 ndint_x_5000_3000 ndint_x_6000_3000 ndint_y_5000_3000 ndint_y_5000_4000 ndint_xy_5000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_6 ndint_x_6000_3000 ndint_x_7000_3000 ndint_y_6000_3000 ndint_y_6000_4000 ndint_xy_6000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_7 ndint_x_7000_3000 ndint_x_8000_3000 ndint_y_7000_3000 ndint_y_7000_4000 ndint_xy_7000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_3_8 ndint_x_8000_3000 ndint_x_9000_3000 ndint_y_8000_3000 ndint_y_8000_4000 ndint_xy_8000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_0 ndint_x_0_4000 ndint_x_1000_4000 ndint_y_0_4000 ndint_y_0_5000 ndint_xy_0_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_1 ndint_x_1000_4000 ndint_x_2000_4000 ndint_y_1000_4000 ndint_y_1000_5000 ndint_xy_1000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_2 ndint_x_2000_4000 ndint_x_3000_4000 ndint_y_2000_4000 ndint_y_2000_5000 ndint_xy_2000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_3 ndint_x_3000_4000 ndint_x_4000_4000 ndint_y_3000_4000 ndint_y_3000_5000 ndint_xy_3000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_4 ndint_x_4000_4000 ndint_x_5000_4000 ndint_y_4000_4000 ndint_y_4000_5000 ndint_xy_4000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_5 ndint_x_5000_4000 ndint_x_6000_4000 ndint_y_5000_4000 ndint_y_5000_5000 ndint_xy_5000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_6 ndint_x_6000_4000 ndint_x_7000_4000 ndint_y_6000_4000 ndint_y_6000_5000 ndint_xy_6000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_7 ndint_x_7000_4000 ndint_x_8000_4000 ndint_y_7000_4000 ndint_y_7000_5000 ndint_xy_7000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_4_8 ndint_x_8000_4000 ndint_x_9000_4000 ndint_y_8000_4000 ndint_y_8000_5000 ndint_xy_8000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_0 ndint_x_0_5000 ndint_x_1000_5000 ndint_y_0_5000 ndint_y_0_6000 ndint_xy_0_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_1 ndint_x_1000_5000 ndint_x_2000_5000 ndint_y_1000_5000 ndint_y_1000_6000 ndint_xy_1000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_2 ndint_x_2000_5000 ndint_x_3000_5000 ndint_y_2000_5000 ndint_y_2000_6000 ndint_xy_2000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_3 ndint_x_3000_5000 ndint_x_4000_5000 ndint_y_3000_5000 ndint_y_3000_6000 ndint_xy_3000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_4 ndint_x_4000_5000 ndint_x_5000_5000 ndint_y_4000_5000 ndint_y_4000_6000 ndint_xy_4000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_5 ndint_x_5000_5000 ndint_x_6000_5000 ndint_y_5000_5000 ndint_y_5000_6000 ndint_xy_5000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_6 ndint_x_6000_5000 ndint_x_7000_5000 ndint_y_6000_5000 ndint_y_6000_6000 ndint_xy_6000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_7 ndint_x_7000_5000 ndint_x_8000_5000 ndint_y_7000_5000 ndint_y_7000_6000 ndint_xy_7000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_5_8 ndint_x_8000_5000 ndint_x_9000_5000 ndint_y_8000_5000 ndint_y_8000_6000 ndint_xy_8000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_0 ndint_x_0_6000 ndint_x_1000_6000 ndint_y_0_6000 ndint_y_0_7000 ndint_xy_0_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_1 ndint_x_1000_6000 ndint_x_2000_6000 ndint_y_1000_6000 ndint_y_1000_7000 ndint_xy_1000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_2 ndint_x_2000_6000 ndint_x_3000_6000 ndint_y_2000_6000 ndint_y_2000_7000 ndint_xy_2000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_3 ndint_x_3000_6000 ndint_x_4000_6000 ndint_y_3000_6000 ndint_y_3000_7000 ndint_xy_3000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_4 ndint_x_4000_6000 ndint_x_5000_6000 ndint_y_4000_6000 ndint_y_4000_7000 ndint_xy_4000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_5 ndint_x_5000_6000 ndint_x_6000_6000 ndint_y_5000_6000 ndint_y_5000_7000 ndint_xy_5000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_6 ndint_x_6000_6000 ndint_x_7000_6000 ndint_y_6000_6000 ndint_y_6000_7000 ndint_xy_6000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_7 ndint_x_7000_6000 ndint_x_8000_6000 ndint_y_7000_6000 ndint_y_7000_7000 ndint_xy_7000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_6_8 ndint_x_8000_6000 ndint_x_9000_6000 ndint_y_8000_6000 ndint_y_8000_7000 ndint_xy_8000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_0 ndint_x_0_7000 ndint_x_1000_7000 ndint_y_0_7000 ndint_y_0_8000 ndint_xy_0_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_1 ndint_x_1000_7000 ndint_x_2000_7000 ndint_y_1000_7000 ndint_y_1000_8000 ndint_xy_1000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_2 ndint_x_2000_7000 ndint_x_3000_7000 ndint_y_2000_7000 ndint_y_2000_8000 ndint_xy_2000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_3 ndint_x_3000_7000 ndint_x_4000_7000 ndint_y_3000_7000 ndint_y_3000_8000 ndint_xy_3000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_4 ndint_x_4000_7000 ndint_x_5000_7000 ndint_y_4000_7000 ndint_y_4000_8000 ndint_xy_4000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_5 ndint_x_5000_7000 ndint_x_6000_7000 ndint_y_5000_7000 ndint_y_5000_8000 ndint_xy_5000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_6 ndint_x_6000_7000 ndint_x_7000_7000 ndint_y_6000_7000 ndint_y_6000_8000 ndint_xy_6000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_7 ndint_x_7000_7000 ndint_x_8000_7000 ndint_y_7000_7000 ndint_y_7000_8000 ndint_xy_7000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_7_8 ndint_x_8000_7000 ndint_x_9000_7000 ndint_y_8000_7000 ndint_y_8000_8000 ndint_xy_8000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_0 ndint_x_0_8000 ndint_x_1000_8000 ndint_y_0_8000 ndint_y_0_9000 ndint_xy_0_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_1 ndint_x_1000_8000 ndint_x_2000_8000 ndint_y_1000_8000 ndint_y_1000_9000 ndint_xy_1000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_2 ndint_x_2000_8000 ndint_x_3000_8000 ndint_y_2000_8000 ndint_y_2000_9000 ndint_xy_2000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_3 ndint_x_3000_8000 ndint_x_4000_8000 ndint_y_3000_8000 ndint_y_3000_9000 ndint_xy_3000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_4 ndint_x_4000_8000 ndint_x_5000_8000 ndint_y_4000_8000 ndint_y_4000_9000 ndint_xy_4000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_5 ndint_x_5000_8000 ndint_x_6000_8000 ndint_y_5000_8000 ndint_y_5000_9000 ndint_xy_5000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_6 ndint_x_6000_8000 ndint_x_7000_8000 ndint_y_6000_8000 ndint_y_6000_9000 ndint_xy_6000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_7 ndint_x_7000_8000 ndint_x_8000_8000 ndint_y_7000_8000 ndint_y_7000_9000 ndint_xy_7000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xdint_8_8 ndint_x_8000_8000 ndint_x_9000_8000 ndint_y_8000_8000 ndint_y_8000_9000 ndint_xy_8000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'

xsint_0_0 nsint_x_0_0 nsint_x_1000_0 nsint_y_0_0 nsint_y_0_1000 nsint_xy_0_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_1 nsint_x_1000_0 nsint_x_2000_0 nsint_y_1000_0 nsint_y_1000_1000 nsint_xy_1000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_2 nsint_x_2000_0 nsint_x_3000_0 nsint_y_2000_0 nsint_y_2000_1000 nsint_xy_2000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_3 nsint_x_3000_0 nsint_x_4000_0 nsint_y_3000_0 nsint_y_3000_1000 nsint_xy_3000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_4 nsint_x_4000_0 nsint_x_5000_0 nsint_y_4000_0 nsint_y_4000_1000 nsint_xy_4000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_5 nsint_x_5000_0 nsint_x_6000_0 nsint_y_5000_0 nsint_y_5000_1000 nsint_xy_5000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_6 nsint_x_6000_0 nsint_x_7000_0 nsint_y_6000_0 nsint_y_6000_1000 nsint_xy_6000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_7 nsint_x_7000_0 nsint_x_8000_0 nsint_y_7000_0 nsint_y_7000_1000 nsint_xy_7000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_0_8 nsint_x_8000_0 nsint_x_9000_0 nsint_y_8000_0 nsint_y_8000_1000 nsint_xy_8000_0 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_0 nsint_x_0_1000 nsint_x_1000_1000 nsint_y_0_1000 nsint_y_0_2000 nsint_xy_0_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_1 nsint_x_1000_1000 nsint_x_2000_1000 nsint_y_1000_1000 nsint_y_1000_2000 nsint_xy_1000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_2 nsint_x_2000_1000 nsint_x_3000_1000 nsint_y_2000_1000 nsint_y_2000_2000 nsint_xy_2000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_3 nsint_x_3000_1000 nsint_x_4000_1000 nsint_y_3000_1000 nsint_y_3000_2000 nsint_xy_3000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_4 nsint_x_4000_1000 nsint_x_5000_1000 nsint_y_4000_1000 nsint_y_4000_2000 nsint_xy_4000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_5 nsint_x_5000_1000 nsint_x_6000_1000 nsint_y_5000_1000 nsint_y_5000_2000 nsint_xy_5000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_6 nsint_x_6000_1000 nsint_x_7000_1000 nsint_y_6000_1000 nsint_y_6000_2000 nsint_xy_6000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_7 nsint_x_7000_1000 nsint_x_8000_1000 nsint_y_7000_1000 nsint_y_7000_2000 nsint_xy_7000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_1_8 nsint_x_8000_1000 nsint_x_9000_1000 nsint_y_8000_1000 nsint_y_8000_2000 nsint_xy_8000_1000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_0 nsint_x_0_2000 nsint_x_1000_2000 nsint_y_0_2000 nsint_y_0_3000 nsint_xy_0_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_1 nsint_x_1000_2000 nsint_x_2000_2000 nsint_y_1000_2000 nsint_y_1000_3000 nsint_xy_1000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_2 nsint_x_2000_2000 nsint_x_3000_2000 nsint_y_2000_2000 nsint_y_2000_3000 nsint_xy_2000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_3 nsint_x_3000_2000 nsint_x_4000_2000 nsint_y_3000_2000 nsint_y_3000_3000 nsint_xy_3000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_4 nsint_x_4000_2000 nsint_x_5000_2000 nsint_y_4000_2000 nsint_y_4000_3000 nsint_xy_4000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_5 nsint_x_5000_2000 nsint_x_6000_2000 nsint_y_5000_2000 nsint_y_5000_3000 nsint_xy_5000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_6 nsint_x_6000_2000 nsint_x_7000_2000 nsint_y_6000_2000 nsint_y_6000_3000 nsint_xy_6000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_7 nsint_x_7000_2000 nsint_x_8000_2000 nsint_y_7000_2000 nsint_y_7000_3000 nsint_xy_7000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_2_8 nsint_x_8000_2000 nsint_x_9000_2000 nsint_y_8000_2000 nsint_y_8000_3000 nsint_xy_8000_2000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_0 nsint_x_0_3000 nsint_x_1000_3000 nsint_y_0_3000 nsint_y_0_4000 nsint_xy_0_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_1 nsint_x_1000_3000 nsint_x_2000_3000 nsint_y_1000_3000 nsint_y_1000_4000 nsint_xy_1000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_2 nsint_x_2000_3000 nsint_x_3000_3000 nsint_y_2000_3000 nsint_y_2000_4000 nsint_xy_2000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_3 nsint_x_3000_3000 nsint_x_4000_3000 nsint_y_3000_3000 nsint_y_3000_4000 nsint_xy_3000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_4 nsint_x_4000_3000 nsint_x_5000_3000 nsint_y_4000_3000 nsint_y_4000_4000 nsint_xy_4000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_5 nsint_x_5000_3000 nsint_x_6000_3000 nsint_y_5000_3000 nsint_y_5000_4000 nsint_xy_5000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_6 nsint_x_6000_3000 nsint_x_7000_3000 nsint_y_6000_3000 nsint_y_6000_4000 nsint_xy_6000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_7 nsint_x_7000_3000 nsint_x_8000_3000 nsint_y_7000_3000 nsint_y_7000_4000 nsint_xy_7000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_3_8 nsint_x_8000_3000 nsint_x_9000_3000 nsint_y_8000_3000 nsint_y_8000_4000 nsint_xy_8000_3000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_0 nsint_x_0_4000 nsint_x_1000_4000 nsint_y_0_4000 nsint_y_0_5000 nsint_xy_0_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_1 nsint_x_1000_4000 nsint_x_2000_4000 nsint_y_1000_4000 nsint_y_1000_5000 nsint_xy_1000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_2 nsint_x_2000_4000 nsint_x_3000_4000 nsint_y_2000_4000 nsint_y_2000_5000 nsint_xy_2000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_3 nsint_x_3000_4000 nsint_x_4000_4000 nsint_y_3000_4000 nsint_y_3000_5000 nsint_xy_3000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_4 nsint_x_4000_4000 nsint_x_5000_4000 nsint_y_4000_4000 nsint_y_4000_5000 nsint_xy_4000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_5 nsint_x_5000_4000 nsint_x_6000_4000 nsint_y_5000_4000 nsint_y_5000_5000 nsint_xy_5000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_6 nsint_x_6000_4000 nsint_x_7000_4000 nsint_y_6000_4000 nsint_y_6000_5000 nsint_xy_6000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_7 nsint_x_7000_4000 nsint_x_8000_4000 nsint_y_7000_4000 nsint_y_7000_5000 nsint_xy_7000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_4_8 nsint_x_8000_4000 nsint_x_9000_4000 nsint_y_8000_4000 nsint_y_8000_5000 nsint_xy_8000_4000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_0 nsint_x_0_5000 nsint_x_1000_5000 nsint_y_0_5000 nsint_y_0_6000 nsint_xy_0_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_1 nsint_x_1000_5000 nsint_x_2000_5000 nsint_y_1000_5000 nsint_y_1000_6000 nsint_xy_1000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_2 nsint_x_2000_5000 nsint_x_3000_5000 nsint_y_2000_5000 nsint_y_2000_6000 nsint_xy_2000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_3 nsint_x_3000_5000 nsint_x_4000_5000 nsint_y_3000_5000 nsint_y_3000_6000 nsint_xy_3000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_4 nsint_x_4000_5000 nsint_x_5000_5000 nsint_y_4000_5000 nsint_y_4000_6000 nsint_xy_4000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_5 nsint_x_5000_5000 nsint_x_6000_5000 nsint_y_5000_5000 nsint_y_5000_6000 nsint_xy_5000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_6 nsint_x_6000_5000 nsint_x_7000_5000 nsint_y_6000_5000 nsint_y_6000_6000 nsint_xy_6000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_7 nsint_x_7000_5000 nsint_x_8000_5000 nsint_y_7000_5000 nsint_y_7000_6000 nsint_xy_7000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_5_8 nsint_x_8000_5000 nsint_x_9000_5000 nsint_y_8000_5000 nsint_y_8000_6000 nsint_xy_8000_5000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_0 nsint_x_0_6000 nsint_x_1000_6000 nsint_y_0_6000 nsint_y_0_7000 nsint_xy_0_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_1 nsint_x_1000_6000 nsint_x_2000_6000 nsint_y_1000_6000 nsint_y_1000_7000 nsint_xy_1000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_2 nsint_x_2000_6000 nsint_x_3000_6000 nsint_y_2000_6000 nsint_y_2000_7000 nsint_xy_2000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_3 nsint_x_3000_6000 nsint_x_4000_6000 nsint_y_3000_6000 nsint_y_3000_7000 nsint_xy_3000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_4 nsint_x_4000_6000 nsint_x_5000_6000 nsint_y_4000_6000 nsint_y_4000_7000 nsint_xy_4000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_5 nsint_x_5000_6000 nsint_x_6000_6000 nsint_y_5000_6000 nsint_y_5000_7000 nsint_xy_5000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_6 nsint_x_6000_6000 nsint_x_7000_6000 nsint_y_6000_6000 nsint_y_6000_7000 nsint_xy_6000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_7 nsint_x_7000_6000 nsint_x_8000_6000 nsint_y_7000_6000 nsint_y_7000_7000 nsint_xy_7000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_6_8 nsint_x_8000_6000 nsint_x_9000_6000 nsint_y_8000_6000 nsint_y_8000_7000 nsint_xy_8000_6000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_0 nsint_x_0_7000 nsint_x_1000_7000 nsint_y_0_7000 nsint_y_0_8000 nsint_xy_0_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_1 nsint_x_1000_7000 nsint_x_2000_7000 nsint_y_1000_7000 nsint_y_1000_8000 nsint_xy_1000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_2 nsint_x_2000_7000 nsint_x_3000_7000 nsint_y_2000_7000 nsint_y_2000_8000 nsint_xy_2000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_3 nsint_x_3000_7000 nsint_x_4000_7000 nsint_y_3000_7000 nsint_y_3000_8000 nsint_xy_3000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_4 nsint_x_4000_7000 nsint_x_5000_7000 nsint_y_4000_7000 nsint_y_4000_8000 nsint_xy_4000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_5 nsint_x_5000_7000 nsint_x_6000_7000 nsint_y_5000_7000 nsint_y_5000_8000 nsint_xy_5000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_6 nsint_x_6000_7000 nsint_x_7000_7000 nsint_y_6000_7000 nsint_y_6000_8000 nsint_xy_6000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_7 nsint_x_7000_7000 nsint_x_8000_7000 nsint_y_7000_7000 nsint_y_7000_8000 nsint_xy_7000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_7_8 nsint_x_8000_7000 nsint_x_9000_7000 nsint_y_8000_7000 nsint_y_8000_8000 nsint_xy_8000_7000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_0 nsint_x_0_8000 nsint_x_1000_8000 nsint_y_0_8000 nsint_y_0_9000 nsint_xy_0_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_1 nsint_x_1000_8000 nsint_x_2000_8000 nsint_y_1000_8000 nsint_y_1000_9000 nsint_xy_1000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_2 nsint_x_2000_8000 nsint_x_3000_8000 nsint_y_2000_8000 nsint_y_2000_9000 nsint_xy_2000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_3 nsint_x_3000_8000 nsint_x_4000_8000 nsint_y_3000_8000 nsint_y_3000_9000 nsint_xy_3000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_4 nsint_x_4000_8000 nsint_x_5000_8000 nsint_y_4000_8000 nsint_y_4000_9000 nsint_xy_4000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_5 nsint_x_5000_8000 nsint_x_6000_8000 nsint_y_5000_8000 nsint_y_5000_9000 nsint_xy_5000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_6 nsint_x_6000_8000 nsint_x_7000_8000 nsint_y_6000_8000 nsint_y_6000_9000 nsint_xy_6000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_7 nsint_x_7000_8000 nsint_x_8000_8000 nsint_y_7000_8000 nsint_y_7000_9000 nsint_xy_7000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'
xsint_8_8 nsint_x_8000_8000 nsint_x_9000_8000 nsint_y_8000_8000 nsint_y_8000_9000 nsint_xy_8000_8000 int_unitcell rval='r_int_cell' lval='l_int_cell' cval='c_int_cell'

.include 'unitcell.subckt'

rs_ubump2via_0_0 ns_chiplet1_pad_0_0 nsint_xy_4000_4000 0.001
rd_ubump2via_0_1 nd_chiplet1_pad_0_1 ndint_y_4000_4000 0.001
rs_ubump2via_0_2 ns_chiplet1_pad_0_2 nsint_y_4000_4000 0.001
rd_ubump2via_0_3 nd_chiplet1_pad_0_3 ndint_y_4000_5000 0.001
rs_ubump2via_0_4 ns_chiplet1_pad_0_4 nsint_y_4000_5000 0.001
rd_ubump2via_0_5 nd_chiplet1_pad_0_5 ndint_y_4000_5000 0.001
rs_ubump2via_0_6 ns_chiplet1_pad_0_6 nsint_y_4000_5000 0.001
rd_ubump2via_0_7 nd_chiplet1_pad_0_7 ndint_y_4000_6000 0.001
rs_ubump2via_0_8 ns_chiplet1_pad_0_8 nsint_y_4000_6000 0.001
rd_ubump2via_0_9 nd_chiplet1_pad_0_9 ndint_y_4000_6000 0.001
rd_ubump2via_1_0 nd_chiplet1_pad_1_0 ndint_y_4000_4000 0.001
rs_ubump2via_1_1 ns_chiplet1_pad_1_1 nsint_xy_4000_4000 0.001
rd_ubump2via_1_2 nd_chiplet1_pad_1_2 ndint_y_4000_4000 0.001
rs_ubump2via_1_3 ns_chiplet1_pad_1_3 nsint_y_4000_5000 0.001
rd_ubump2via_1_4 nd_chiplet1_pad_1_4 ndint_y_4000_5000 0.001
rs_ubump2via_1_5 ns_chiplet1_pad_1_5 nsint_y_4000_5000 0.001
rd_ubump2via_1_6 nd_chiplet1_pad_1_6 ndint_y_4000_5000 0.001
rs_ubump2via_1_7 ns_chiplet1_pad_1_7 nsint_y_4000_6000 0.001
rd_ubump2via_1_8 nd_chiplet1_pad_1_8 ndint_y_4000_6000 0.001
rs_ubump2via_1_9 ns_chiplet1_pad_1_9 nsint_y_4000_6000 0.001
rs_ubump2via_2_0 ns_chiplet1_pad_2_0 nsint_y_4000_4000 0.001
rd_ubump2via_2_1 nd_chiplet1_pad_2_1 ndint_y_4000_4000 0.001
rs_ubump2via_2_2 ns_chiplet1_pad_2_2 nsint_xy_4000_4000 0.001
rd_ubump2via_2_3 nd_chiplet1_pad_2_3 ndint_y_4000_5000 0.001
rs_ubump2via_2_4 ns_chiplet1_pad_2_4 nsint_y_4000_5000 0.001
rd_ubump2via_2_5 nd_chiplet1_pad_2_5 ndint_y_4000_5000 0.001
rs_ubump2via_2_6 ns_chiplet1_pad_2_6 nsint_y_4000_5000 0.001
rd_ubump2via_2_7 nd_chiplet1_pad_2_7 ndint_y_4000_6000 0.001
rs_ubump2via_2_8 ns_chiplet1_pad_2_8 nsint_y_4000_6000 0.001
rd_ubump2via_2_9 nd_chiplet1_pad_2_9 ndint_y_4000_6000 0.001
rd_ubump2via_3_0 nd_chiplet1_pad_3_0 ndint_y_5000_4000 0.001
rs_ubump2via_3_1 ns_chiplet1_pad_3_1 nsint_y_5000_4000 0.001
rd_ubump2via_3_2 nd_chiplet1_pad_3_2 ndint_y_5000_4000 0.001
rs_ubump2via_3_3 ns_chiplet1_pad_3_3 nsint_xy_5000_5000 0.001
rd_ubump2via_3_4 nd_chiplet1_pad_3_4 ndint_y_5000_5000 0.001
rs_ubump2via_3_5 ns_chiplet1_pad_3_5 nsint_y_5000_5000 0.001
rd_ubump2via_3_6 nd_chiplet1_pad_3_6 ndint_y_5000_5000 0.001
rs_ubump2via_3_7 ns_chiplet1_pad_3_7 nsint_y_5000_6000 0.001
rd_ubump2via_3_8 nd_chiplet1_pad_3_8 ndint_y_5000_6000 0.001
rs_ubump2via_3_9 ns_chiplet1_pad_3_9 nsint_y_5000_6000 0.001
rs_ubump2via_4_0 ns_chiplet1_pad_4_0 nsint_y_5000_4000 0.001
rd_ubump2via_4_1 nd_chiplet1_pad_4_1 ndint_y_5000_4000 0.001
rs_ubump2via_4_2 ns_chiplet1_pad_4_2 nsint_y_5000_4000 0.001
rd_ubump2via_4_3 nd_chiplet1_pad_4_3 ndint_y_5000_5000 0.001
rs_ubump2via_4_4 ns_chiplet1_pad_4_4 nsint_xy_5000_5000 0.001
rd_ubump2via_4_5 nd_chiplet1_pad_4_5 ndint_y_5000_5000 0.001
rs_ubump2via_4_6 ns_chiplet1_pad_4_6 nsint_y_5000_5000 0.001
rd_ubump2via_4_7 nd_chiplet1_pad_4_7 ndint_y_5000_6000 0.001
rs_ubump2via_4_8 ns_chiplet1_pad_4_8 nsint_y_5000_6000 0.001
rd_ubump2via_4_9 nd_chiplet1_pad_4_9 ndint_y_5000_6000 0.001
rd_ubump2via_5_0 nd_chiplet1_pad_5_0 ndint_y_5000_4000 0.001
rs_ubump2via_5_1 ns_chiplet1_pad_5_1 nsint_y_5000_4000 0.001
rd_ubump2via_5_2 nd_chiplet1_pad_5_2 ndint_y_5000_4000 0.001
rs_ubump2via_5_3 ns_chiplet1_pad_5_3 nsint_y_5000_5000 0.001
rd_ubump2via_5_4 nd_chiplet1_pad_5_4 ndint_y_5000_5000 0.001
rs_ubump2via_5_5 ns_chiplet1_pad_5_5 nsint_xy_5000_5000 0.001
rd_ubump2via_5_6 nd_chiplet1_pad_5_6 ndint_y_5000_5000 0.001
rs_ubump2via_5_7 ns_chiplet1_pad_5_7 nsint_y_5000_6000 0.001
rd_ubump2via_5_8 nd_chiplet1_pad_5_8 ndint_y_5000_6000 0.001
rs_ubump2via_5_9 ns_chiplet1_pad_5_9 nsint_y_5000_6000 0.001
rs_ubump2via_6_0 ns_chiplet1_pad_6_0 nsint_y_5000_4000 0.001
rd_ubump2via_6_1 nd_chiplet1_pad_6_1 ndint_y_5000_4000 0.001
rs_ubump2via_6_2 ns_chiplet1_pad_6_2 nsint_y_5000_4000 0.001
rd_ubump2via_6_3 nd_chiplet1_pad_6_3 ndint_y_5000_5000 0.001
rs_ubump2via_6_4 ns_chiplet1_pad_6_4 nsint_y_5000_5000 0.001
rd_ubump2via_6_5 nd_chiplet1_pad_6_5 ndint_y_5000_5000 0.001
rs_ubump2via_6_6 ns_chiplet1_pad_6_6 nsint_xy_5000_5000 0.001
rd_ubump2via_6_7 nd_chiplet1_pad_6_7 ndint_y_5000_6000 0.001
rs_ubump2via_6_8 ns_chiplet1_pad_6_8 nsint_y_5000_6000 0.001
rd_ubump2via_6_9 nd_chiplet1_pad_6_9 ndint_y_5000_6000 0.001
rd_ubump2via_7_0 nd_chiplet1_pad_7_0 ndint_y_6000_4000 0.001
rs_ubump2via_7_1 ns_chiplet1_pad_7_1 nsint_y_6000_4000 0.001
rd_ubump2via_7_2 nd_chiplet1_pad_7_2 ndint_y_6000_4000 0.001
rs_ubump2via_7_3 ns_chiplet1_pad_7_3 nsint_y_6000_5000 0.001
rd_ubump2via_7_4 nd_chiplet1_pad_7_4 ndint_y_6000_5000 0.001
rs_ubump2via_7_5 ns_chiplet1_pad_7_5 nsint_y_6000_5000 0.001
rd_ubump2via_7_6 nd_chiplet1_pad_7_6 ndint_y_6000_5000 0.001
rs_ubump2via_7_7 ns_chiplet1_pad_7_7 nsint_xy_6000_6000 0.001
rd_ubump2via_7_8 nd_chiplet1_pad_7_8 ndint_y_6000_6000 0.001
rs_ubump2via_7_9 ns_chiplet1_pad_7_9 nsint_y_6000_6000 0.001
rs_ubump2via_8_0 ns_chiplet1_pad_8_0 nsint_y_6000_4000 0.001
rd_ubump2via_8_1 nd_chiplet1_pad_8_1 ndint_y_6000_4000 0.001
rs_ubump2via_8_2 ns_chiplet1_pad_8_2 nsint_y_6000_4000 0.001
rd_ubump2via_8_3 nd_chiplet1_pad_8_3 ndint_y_6000_5000 0.001
rs_ubump2via_8_4 ns_chiplet1_pad_8_4 nsint_y_6000_5000 0.001
rd_ubump2via_8_5 nd_chiplet1_pad_8_5 ndint_y_6000_5000 0.001
rs_ubump2via_8_6 ns_chiplet1_pad_8_6 nsint_y_6000_5000 0.001
rd_ubump2via_8_7 nd_chiplet1_pad_8_7 ndint_y_6000_6000 0.001
rs_ubump2via_8_8 ns_chiplet1_pad_8_8 nsint_xy_6000_6000 0.001
rd_ubump2via_8_9 nd_chiplet1_pad_8_9 ndint_y_6000_6000 0.001
rd_ubump2via_9_0 nd_chiplet1_pad_9_0 ndint_y_6000_4000 0.001
rs_ubump2via_9_1 ns_chiplet1_pad_9_1 nsint_y_6000_4000 0.001
rd_ubump2via_9_2 nd_chiplet1_pad_9_2 ndint_y_6000_4000 0.001
rs_ubump2via_9_3 ns_chiplet1_pad_9_3 nsint_y_6000_5000 0.001
rd_ubump2via_9_4 nd_chiplet1_pad_9_4 ndint_y_6000_5000 0.001
rs_ubump2via_9_5 ns_chiplet1_pad_9_5 nsint_y_6000_5000 0.001
rd_ubump2via_9_6 nd_chiplet1_pad_9_6 ndint_y_6000_5000 0.001
rs_ubump2via_9_7 ns_chiplet1_pad_9_7 nsint_y_6000_6000 0.001
rd_ubump2via_9_8 nd_chiplet1_pad_9_8 ndint_y_6000_6000 0.001
rs_ubump2via_9_9 ns_chiplet1_pad_9_9 nsint_xy_6000_6000 0.001

*-- chiplet instance [0]: chiplet1
xchiplet_chiplet1
+ns_chiplet1_pad_0_0
+nd_chiplet1_pad_0_1
+ns_chiplet1_pad_0_2
+nd_chiplet1_pad_0_3
+ns_chiplet1_pad_0_4
+nd_chiplet1_pad_0_5
+ns_chiplet1_pad_0_6
+nd_chiplet1_pad_0_7
+ns_chiplet1_pad_0_8
+nd_chiplet1_pad_0_9
+nd_chiplet1_pad_1_0
+ns_chiplet1_pad_1_1
+nd_chiplet1_pad_1_2
+ns_chiplet1_pad_1_3
+nd_chiplet1_pad_1_4
+ns_chiplet1_pad_1_5
+nd_chiplet1_pad_1_6
+ns_chiplet1_pad_1_7
+nd_chiplet1_pad_1_8
+ns_chiplet1_pad_1_9
+ns_chiplet1_pad_2_0
+nd_chiplet1_pad_2_1
+ns_chiplet1_pad_2_2
+nd_chiplet1_pad_2_3
+ns_chiplet1_pad_2_4
+nd_chiplet1_pad_2_5
+ns_chiplet1_pad_2_6
+nd_chiplet1_pad_2_7
+ns_chiplet1_pad_2_8
+nd_chiplet1_pad_2_9
+nd_chiplet1_pad_3_0
+ns_chiplet1_pad_3_1
+nd_chiplet1_pad_3_2
+ns_chiplet1_pad_3_3
+nd_chiplet1_pad_3_4
+ns_chiplet1_pad_3_5
+nd_chiplet1_pad_3_6
+ns_chiplet1_pad_3_7
+nd_chiplet1_pad_3_8
+ns_chiplet1_pad_3_9
+ns_chiplet1_pad_4_0
+nd_chiplet1_pad_4_1
+ns_chiplet1_pad_4_2
+nd_chiplet1_pad_4_3
+ns_chiplet1_pad_4_4
+nd_chiplet1_pad_4_5
+ns_chiplet1_pad_4_6
+nd_chiplet1_pad_4_7
+ns_chiplet1_pad_4_8
+nd_chiplet1_pad_4_9
+nd_chiplet1_pad_5_0
+ns_chiplet1_pad_5_1
+nd_chiplet1_pad_5_2
+ns_chiplet1_pad_5_3
+nd_chiplet1_pad_5_4
+ns_chiplet1_pad_5_5
+nd_chiplet1_pad_5_6
+ns_chiplet1_pad_5_7
+nd_chiplet1_pad_5_8
+ns_chiplet1_pad_5_9
+ns_chiplet1_pad_6_0
+nd_chiplet1_pad_6_1
+ns_chiplet1_pad_6_2
+nd_chiplet1_pad_6_3
+ns_chiplet1_pad_6_4
+nd_chiplet1_pad_6_5
+ns_chiplet1_pad_6_6
+nd_chiplet1_pad_6_7
+ns_chiplet1_pad_6_8
+nd_chiplet1_pad_6_9
+nd_chiplet1_pad_7_0
+ns_chiplet1_pad_7_1
+nd_chiplet1_pad_7_2
+ns_chiplet1_pad_7_3
+nd_chiplet1_pad_7_4
+ns_chiplet1_pad_7_5
+nd_chiplet1_pad_7_6
+ns_chiplet1_pad_7_7
+nd_chiplet1_pad_7_8
+ns_chiplet1_pad_7_9
+ns_chiplet1_pad_8_0
+nd_chiplet1_pad_8_1
+ns_chiplet1_pad_8_2
+nd_chiplet1_pad_8_3
+ns_chiplet1_pad_8_4
+nd_chiplet1_pad_8_5
+ns_chiplet1_pad_8_6
+nd_chiplet1_pad_8_7
+ns_chiplet1_pad_8_8
+nd_chiplet1_pad_8_9
+nd_chiplet1_pad_9_0
+ns_chiplet1_pad_9_1
+nd_chiplet1_pad_9_2
+ns_chiplet1_pad_9_3
+nd_chiplet1_pad_9_4
+ns_chiplet1_pad_9_5
+nd_chiplet1_pad_9_6
+ns_chiplet1_pad_9_7
+nd_chiplet1_pad_9_8
+ns_chiplet1_pad_9_9
+chiplet1
.include 'chiplet1_ac.subckt'

*-- tsv array
xsint_tsv_0_0 nsint_tsv_0_0 nsint_bump_0_0 int_tsv
xdint_tsv_0_1 ndint_tsv_0_1 ndint_bump_0_1 int_tsv
xsint_tsv_0_2 nsint_tsv_0_2 nsint_bump_0_2 int_tsv
xdint_tsv_0_3 ndint_tsv_0_3 ndint_bump_0_3 int_tsv
xsint_tsv_0_4 nsint_tsv_0_4 nsint_bump_0_4 int_tsv
xdint_tsv_1_0 ndint_tsv_1_0 ndint_bump_1_0 int_tsv
xsint_tsv_1_1 nsint_tsv_1_1 nsint_bump_1_1 int_tsv
xdint_tsv_1_2 ndint_tsv_1_2 ndint_bump_1_2 int_tsv
xsint_tsv_1_3 nsint_tsv_1_3 nsint_bump_1_3 int_tsv
xdint_tsv_1_4 ndint_tsv_1_4 ndint_bump_1_4 int_tsv
xsint_tsv_2_0 nsint_tsv_2_0 nsint_bump_2_0 int_tsv
xdint_tsv_2_1 ndint_tsv_2_1 ndint_bump_2_1 int_tsv
xsint_tsv_2_2 nsint_tsv_2_2 nsint_bump_2_2 int_tsv
xdint_tsv_2_3 ndint_tsv_2_3 ndint_bump_2_3 int_tsv
xsint_tsv_2_4 nsint_tsv_2_4 nsint_bump_2_4 int_tsv
xdint_tsv_3_0 ndint_tsv_3_0 ndint_bump_3_0 int_tsv
xsint_tsv_3_1 nsint_tsv_3_1 nsint_bump_3_1 int_tsv
xdint_tsv_3_2 ndint_tsv_3_2 ndint_bump_3_2 int_tsv
xsint_tsv_3_3 nsint_tsv_3_3 nsint_bump_3_3 int_tsv
xdint_tsv_3_4 ndint_tsv_3_4 ndint_bump_3_4 int_tsv
xsint_tsv_4_0 nsint_tsv_4_0 nsint_bump_4_0 int_tsv
xdint_tsv_4_1 ndint_tsv_4_1 ndint_bump_4_1 int_tsv
xsint_tsv_4_2 nsint_tsv_4_2 nsint_bump_4_2 int_tsv
xdint_tsv_4_3 ndint_tsv_4_3 ndint_bump_4_3 int_tsv
xsint_tsv_4_4 nsint_tsv_4_4 nsint_bump_4_4 int_tsv
.include 'int_tsv.subckt'

*-- tsv to via
rsint_tsv2via_0_0 nsint_tsv_0_0 nsint_xy_2000_2000 0.001
rdint_tsv2via_0_1 ndint_tsv_0_1 ndint_y_2000_3000 0.001
rsint_tsv2via_0_2 nsint_tsv_0_2 nsint_y_2000_5000 0.001
rdint_tsv2via_0_3 ndint_tsv_0_3 ndint_xy_2000_7000 0.001
rsint_tsv2via_0_4 nsint_tsv_0_4 nsint_y_2000_8000 0.001
rdint_tsv2via_1_0 ndint_tsv_1_0 ndint_y_3000_2000 0.001
rsint_tsv2via_1_1 nsint_tsv_1_1 nsint_xy_3000_3000 0.001
rdint_tsv2via_1_2 ndint_tsv_1_2 ndint_y_3000_5000 0.001
rsint_tsv2via_1_3 nsint_tsv_1_3 nsint_y_3000_7000 0.001
rdint_tsv2via_1_4 ndint_tsv_1_4 ndint_xy_3000_8000 0.001
rsint_tsv2via_2_0 nsint_tsv_2_0 nsint_y_5000_2000 0.001
rdint_tsv2via_2_1 ndint_tsv_2_1 ndint_y_5000_3000 0.001
rsint_tsv2via_2_2 nsint_tsv_2_2 nsint_xy_5000_5000 0.001
rdint_tsv2via_2_3 ndint_tsv_2_3 ndint_y_5000_7000 0.001
rsint_tsv2via_2_4 nsint_tsv_2_4 nsint_y_5000_8000 0.001
rdint_tsv2via_3_0 ndint_tsv_3_0 ndint_xy_7000_2000 0.001
rsint_tsv2via_3_1 nsint_tsv_3_1 nsint_y_7000_3000 0.001
rdint_tsv2via_3_2 ndint_tsv_3_2 ndint_y_7000_5000 0.001
rsint_tsv2via_3_3 nsint_tsv_3_3 nsint_xy_7000_7000 0.001
rdint_tsv2via_3_4 ndint_tsv_3_4 ndint_y_7000_8000 0.001
rsint_tsv2via_4_0 nsint_tsv_4_0 nsint_y_8000_2000 0.001
rdint_tsv2via_4_1 ndint_tsv_4_1 ndint_xy_8000_3000 0.001
rsint_tsv2via_4_2 nsint_tsv_4_2 nsint_y_8000_5000 0.001
rdint_tsv2via_4_3 ndint_tsv_4_3 ndint_y_8000_7000 0.001
rsint_tsv2via_4_4 nsint_tsv_4_4 nsint_xy_8000_8000 0.001

*-- tsv bump array to pkg
rsint_tsv_0_0 nsint_bump_0_0 ns_pkg_pad 0.001
rdint_tsv_0_1 ndint_bump_0_1 nd_pkg_pad 0.001
rsint_tsv_0_2 nsint_bump_0_2 ns_pkg_pad 0.001
rdint_tsv_0_3 ndint_bump_0_3 nd_pkg_pad 0.001
rsint_tsv_0_4 nsint_bump_0_4 ns_pkg_pad 0.001
rdint_tsv_1_0 ndint_bump_1_0 nd_pkg_pad 0.001
rsint_tsv_1_1 nsint_bump_1_1 ns_pkg_pad 0.001
rdint_tsv_1_2 ndint_bump_1_2 nd_pkg_pad 0.001
rsint_tsv_1_3 nsint_bump_1_3 ns_pkg_pad 0.001
rdint_tsv_1_4 ndint_bump_1_4 nd_pkg_pad 0.001
rsint_tsv_2_0 nsint_bump_2_0 ns_pkg_pad 0.001
rdint_tsv_2_1 ndint_bump_2_1 nd_pkg_pad 0.001
rsint_tsv_2_2 nsint_bump_2_2 ns_pkg_pad 0.001
rdint_tsv_2_3 ndint_bump_2_3 nd_pkg_pad 0.001
rsint_tsv_2_4 nsint_bump_2_4 ns_pkg_pad 0.001
rdint_tsv_3_0 ndint_bump_3_0 nd_pkg_pad 0.001
rsint_tsv_3_1 nsint_bump_3_1 ns_pkg_pad 0.001
rdint_tsv_3_2 ndint_bump_3_2 nd_pkg_pad 0.001
rsint_tsv_3_3 nsint_bump_3_3 ns_pkg_pad 0.001
rdint_tsv_3_4 ndint_bump_3_4 nd_pkg_pad 0.001
rsint_tsv_4_0 nsint_bump_4_0 ns_pkg_pad 0.001
rdint_tsv_4_1 ndint_bump_4_1 nd_pkg_pad 0.001
rsint_tsv_4_2 nsint_bump_4_2 ns_pkg_pad 0.001
rdint_tsv_4_3 ndint_bump_4_3 nd_pkg_pad 0.001
rsint_tsv_4_4 nsint_bump_4_4 ns_pkg_pad 0.001

*-- pkg instances
xpkg_vdd vdd_pkg nd_pkg_pad pkg_model
xpkg_vss vss_pkg ns_pkg_pad pkg_model
.include 'pkg.subckt'

*-- pcb instances
xpcb_vdd vdd vdd_pkg pcb_model
xpcb_vss vss vss_pkg pcb_model
.include 'pcb.subckt'


*-- external power source
ivdd 0 vdd 0 ac 1
ivss 0 vss 0 ac 1
.ac dec 100 1e+06 1e+10
.end
